52	24
shingles	yexeyexeyexeyexeyexeyexe	aaxexeyexeyexeyexexexeye	yeyeCeyeCeyeCeyeCeBeCeCe	aaxexeyexeyexeye	CfyfxeoeoeoeCexeCeyeyeCe	yexeyeyexeyexeyeyexeyexe	yexeyexeyexeyexexeyeyexe	xexexeyexeyexeyexeyexexe	yfxeyeyexexeyexeyexexeye	aaxexeyexeqe	CfCfCfCfCeyeCeCeyeCeyeCe	xexeyeyOra	yeyeyera	aayOqe	xeCeyeyeCeCfxeyeyeyfCeye	yexexeyeyexexexexexexexe	aayO	yexexeyexeyexeyexeyexeye	CeoeCfCeCeyfCeyeyeCeCeyf	xexeyeyexeyeyexeyeyexeye	CfxeyeyeyfCeyeCeCeyeCeye	aaqe	xeyexeyeyeyexeyexeyeyeye	aaxexeyexeyexeyexeyexeyf	yeyexeyexeyeyeyexeyexeye	CfCfCfCfCfCfCfCfCfCfCfCf	CfCfCfCeCeyfCfCeCeyeyeCe	xexeyeyeyexeyeyeyeyeyeye	aaCOyOxeyeyeye	aayOCeraHayOCeyO	yeyeCeCeyfCfyfxeoeoeoeCe	CeyfCfyfxeoeoeoeCexeCeye	xeCexexexexexeyeyexeyeye	aaxexeyexeyexeyexeyexeye	xeyeyexexeyeyexexeyeyexe	xeyexeyexexeyexeyexexeye	aaxexeyexexeyexeyexeyexe	xeyeyeyfyfyfyfCexeyeyexe	yexeyexeyexeyexe	xexeyeyeyexeyeyeyeyeyeCe	xeyexexeoeoeoeCexeCeyeye	yeyeCeCeyeCeyeCeCeoeBeCe	CeCeoeBeCeCeoeCfCeCeyfCe	yeyexeyeyeyexeyeyeyeyeye	CeCfxeyeyeyfCeCeCeCeCeCe	oeoeCexeCeyeyeCeCfxeyeye	yeCfyfyeyeCeCeyfCfyfxeoe	yfCfCfCfCfCfCfCfCfCfCfCf	CfCfCfCfCeyeyfyfCfCeCfCf	CeoeBeCeCeoeCfCfCfCfCfCf	yeCeCfyfCeyeCeCeyeCeyeCe	yeCeCeCeoeBeoeCeCeyfxeoe
0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	1	0	0	0	0	0	0	0	0	0	0	0	1	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0
1	0	0	0	0	0	0	0	0	0	0	0	0	0	2	0	0	0	0	0	0	0	1	0	0	0	0	0	0	0	1	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0
2	0	0	0	0	0	1	1	1	0	0	0	0	1	0	0	1	0	1	0	1	0	1	1	0	1	0	0	1	0	0	0	0	1	1	1	2	0	0	0	0	0	0	0	1	0	0	0	0	0	0	0	0
3	0	0	0	0	0	0	0	0	0	1	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0
4	0	0	0	1	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0
5	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	1	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0
6	0	0	1	0	1	0	0	0	1	0	1	0	0	0	1	0	0	0	1	0	1	0	0	1	0	1	1	0	0	0	1	1	0	0	0	0	0	1	0	1	1	1	1	0	1	1	1	1	1	1	1	1
7	0	1	0	0	0	0	0	0	0	0	0	1	0	0	0	0	0	0	0	0	0	1	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0
8	0	0	0	0	0	1	1	1	0	0	0	0	1	0	0	1	0	1	0	1	0	1	1	0	1	0	0	1	0	0	0	0	1	1	1	2	0	0	0	0	0	0	0	1	0	0	0	0	0	0	0	0
9	18	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	0	1	0	1	0	0	0	0	0	0	0	0	0	0	0	0	0
